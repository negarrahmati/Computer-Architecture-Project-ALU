module ICache(address,data_out);
	parameter WIDTH = 32;
	parameter SIZE = 108;
	parameter WIDTH_ADD = 32;
	parameter BYTE = 8;
	
	input [WIDTH_ADD-1:0] address;
	
	output [WIDTH-1:0] data_out;
	
	reg [BYTE-1:0] mem [SIZE-1:0];
	
	assign	data_out = {{mem[address+3]},{mem[address+2]},{mem[address+1]},{mem[address]}};
	
	initial 
	begin
/*		mem[3][BYTE-1:0] = 8'b11100000;
		mem[2][BYTE-1:0] = 8'b00100010;
		mem[1][BYTE-1:0] = 8'b00000000;
		mem[0][BYTE-1:0] = 8'b00001111;
		mem[7][BYTE-1:0] = 8'b11111111;
		mem[6][BYTE-1:0] = 8'b11111111;
		mem[5][BYTE-1:0] = 8'b11111111;
		mem[4][BYTE-1:0] = 8'b11111111;*/

		mem[3][BYTE-1:0] = 8'b11100000;
		mem[2][BYTE-1:0] = 8'b00100001;
		mem[1][BYTE-1:0] = 8'b00000000;
		mem[0][BYTE-1:0] = 8'b00000100;
		mem[7][BYTE-1:0] = 8'b11100000;
		mem[6][BYTE-1:0] = 8'b01000010;
		mem[5][BYTE-1:0] = 8'b00000000;
		mem[4][BYTE-1:0] = 8'b00000101;
		mem[11][BYTE-1:0] = 8'b00000000;
		mem[10][BYTE-1:0] = 8'b00100010;
		mem[9][BYTE-1:0] = 8'b10101000;
		mem[8][BYTE-1:0] = 8'b00000000;
		mem[15][BYTE-1:0] = 8'b00000000;
		mem[14][BYTE-1:0] = 8'b00100010;
		mem[13][BYTE-1:0] = 8'b10110000;
		mem[12][BYTE-1:0] = 8'b00000001;
		mem[19][BYTE-1:0] = 8'b11101000;
		mem[18][BYTE-1:0] = 8'b00010101;
		mem[17][BYTE-1:0] = 8'b00000000;
		mem[16][BYTE-1:0] = 8'b00000000;
		mem[23][BYTE-1:0] = 8'b11101000;
		mem[22][BYTE-1:0] = 8'b00110110;
		mem[21][BYTE-1:0] = 8'b00000000;
		mem[20][BYTE-1:0] = 8'b00000000;
		mem[27][BYTE-1:0] = 8'b11100100;
		mem[26][BYTE-1:0] = 8'b00010111;
		mem[25][BYTE-1:0] = 8'b00000000;
		mem[24][BYTE-1:0] = 8'b00000000;
		mem[31][BYTE-1:0] = 8'b00000010;
		mem[30][BYTE-1:0] = 8'b11100000;
		mem[29][BYTE-1:0] = 8'b10111000;
		mem[28][BYTE-1:0] = 8'b10001100;
		mem[35][BYTE-1:0] = 8'b11101000;
		mem[34][BYTE-1:0] = 8'b00110111;
		mem[33][BYTE-1:0] = 8'b00000000;
		mem[32][BYTE-1:0] = 8'b00000100;
		mem[39][BYTE-1:0] = 8'b00000010;
		mem[38][BYTE-1:0] = 8'b11100000;
		mem[37][BYTE-1:0] = 8'b10111001;
		mem[36][BYTE-1:0] = 8'b00001101;
		mem[43][BYTE-1:0] = 8'b11101000;
		mem[42][BYTE-1:0] = 8'b00110111;
		mem[41][BYTE-1:0] = 8'b00000000;
		mem[40][BYTE-1:0] = 8'b00001000;
		mem[47][BYTE-1:0] = 8'b11100000;
		mem[46][BYTE-1:0] = 8'b01100011;
		mem[45][BYTE-1:0] = 8'b00000000;
		mem[44][BYTE-1:0] = 8'b00100010;
		mem[51][BYTE-1:0] = 8'b11100000;
		mem[50][BYTE-1:0] = 8'b10000100;
		mem[49][BYTE-1:0] = 8'b00000000;
		mem[48][BYTE-1:0] = 8'b00101101;
		mem[55][BYTE-1:0] = 8'b11001100;
		mem[54][BYTE-1:0] = 8'b10000011;
		mem[53][BYTE-1:0] = 8'b00000000;
		mem[52][BYTE-1:0] = 8'b00000010;
		mem[59][BYTE-1:0] = 8'b11101000;
		mem[58][BYTE-1:0] = 8'b00100011;
		mem[57][BYTE-1:0] = 8'b00000000;
		mem[56][BYTE-1:0] = 8'b00001100;
		mem[63][BYTE-1:0] = 8'b10000000;
		mem[62][BYTE-1:0] = 8'b00000000;
		mem[61][BYTE-1:0] = 8'b00000000;
		mem[60][BYTE-1:0] = 8'b00010001;
		mem[67][BYTE-1:0] = 8'b11101000;
		mem[66][BYTE-1:0] = 8'b00100100;
		mem[65][BYTE-1:0] = 8'b00000000;
		mem[64][BYTE-1:0] = 8'b00001100;
		mem[71][BYTE-1:0] = 8'b11010000;
		mem[70][BYTE-1:0] = 8'b01100100;
		mem[69][BYTE-1:0] = 8'b00000000;
		mem[68][BYTE-1:0] = 8'b00000010;
		mem[75][BYTE-1:0] = 8'b11101000;
		mem[74][BYTE-1:0] = 8'b00100011;
		mem[73][BYTE-1:0] = 8'b00000000;
		mem[72][BYTE-1:0] = 8'b00010000;
		mem[79][BYTE-1:0] = 8'b10000000;
		mem[78][BYTE-1:0] = 8'b00000000;
		mem[77][BYTE-1:0] = 8'b00000000;
		mem[76][BYTE-1:0] = 8'b00010101;
		mem[83][BYTE-1:0] = 8'b11101000;
		mem[82][BYTE-1:0] = 8'b00100100;
		mem[81][BYTE-1:0] = 8'b00000000;
		mem[80][BYTE-1:0] = 8'b00010000;
		mem[87][BYTE-1:0] = 8'b10000100;
		mem[86][BYTE-1:0] = 8'b00000000;
		mem[85][BYTE-1:0] = 8'b00000000;
		mem[84][BYTE-1:0] = 8'b00011000;
		mem[91][BYTE-1:0] = 8'b11100000;
		mem[90][BYTE-1:0] = 8'b01100011;
		mem[89][BYTE-1:0] = 8'b00000000;
		mem[88][BYTE-1:0] = 8'b00001011;
		mem[95][BYTE-1:0] = 8'b11101000;
		mem[94][BYTE-1:0] = 8'b00100011;
		mem[93][BYTE-1:0] = 8'b00000000;
		mem[92][BYTE-1:0] = 8'b00010100;
		mem[99][BYTE-1:0] = 8'b11001100;
		mem[98][BYTE-1:0] = 8'b10000011;
		mem[97][BYTE-1:0] = 8'b00000000;
		mem[96][BYTE-1:0] = 8'b00000001;
		mem[103][BYTE-1:0] = 8'b000000_00;
		mem[102][BYTE-1:0] = 8'b000_00000;
		mem[101][BYTE-1:0] = 8'b00000000;
		mem[100][BYTE-1:0] = 8'b0000_1_000;
		mem[107][BYTE-1:0] = 8'b11111111;
		mem[106][BYTE-1:0] = 8'b11111111;
		mem[105][BYTE-1:0] = 8'b11111111;
		mem[104][BYTE-1:0] = 8'b11111111;		
	end
endmodule 